** sch_path: /foss/designs/sky130_ota_5t/xschem/sky130_ota_5t.sch
.subckt sky130_ota_5t Vp Vn Vout VDD VSS Ib
*.PININFO Vp:I Vn:I Vout:O VDD:B VSS:B Ib:I
XM4 net1 Vp node VSS sky130_fd_pr__nfet_01v8 L=0.5 W=20 nf=4 m=1
XM1 Vout net1 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 m=1
XM2 net1 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 m=1
XM3 Vout Vn node VSS sky130_fd_pr__nfet_01v8 L=0.5 W=20 nf=4 m=1
XM5 node Ib VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=2 m=1
XM6 Ib Ib VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=2 m=1
XM7 Vout VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 m=1
XM8 node VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.5 W=20 nf=4 m=1
XM9 node VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=2 m=1
.ends
.end
